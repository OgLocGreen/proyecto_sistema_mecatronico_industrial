PLL_servo_inst : PLL_servo PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
